library verilog;
use verilog.vl_types.all;
entity FINALPROCESSOR_vlg_vec_tst is
end FINALPROCESSOR_vlg_vec_tst;
